`timescale 1ns/1ps



module top();
complex_matrix_hermitian u0();
complex_matrix_multiplier u1();
complex_matrix_multiplier_zeroed u15();
complex_matrix_adder_parallel u2();
scalar_divide u3();
complex_matrix_mult_4_mult u4();

endmodule