`timescale 1ns/1ps



module top();
complex_matrix_multiplier u1();
complex_matrix_multiplier_zeroed u15();
complex_matrix_adder_parallel u2();
scalar_divide_const u3();
scalar_divide u35();
complex_matrix_mult_1_mult u4();
matrix_accumulator_no_latency u5();
rxx u7();
p_theta u8();
bartlett_time_domain u9();


endmodule